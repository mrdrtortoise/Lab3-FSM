module lfsr_7 (
    input   logic       clk,
    input   logic       rst_l,
    input   logic       en,
    output  logic [6:0] data_out
);

logic [6:0] sreg;

always_ff @( posedge clk, posedge rst_l ) begin
    if(rst_l) begin
        sreg <= 7'b1;
    end
    else if(en)begin
        sreg <= {sreg[5:0], sreg[6] ^ sreg[2]};
    end
    
end
assign data_out = sreg;
endmodule
